`define MDF_OP_WIDTH 4
`define MDF_OP_MUL `MDF_OP_WIDTH'd0
`define MDF_OP_DIV `MDF_OP_WIDTH'd1
`define MDF_OP_NOP `MDF_OP_WIDTH'd2
`define MDF_OP_SGN `MDF_OP_WIDTH'd3

`define MD_OUT_LO  1'b0
`define MD_OUT_HI  1'b1

